

module ethernet: 


endmodule